
module detect_22kHz(clk,clk_out);
input clk;
output clk_out;

endmodule 